`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: Evan Nguyen
// 
// Create Date: 11/30/2021 12:32:32 AM
// Design Name: 
// Module Name: game_of_life
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: Open sourced from Spencer Elliot. Revisioned for FPGA implementation for 
//              CSULB's CECS 361 Final Project by Evan Nguyen.
//              Game of life algorithm with presets. 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


/**
 * Main module to be instantiated in a project that uses a VGA controller
 */
module game_of_life(KEY, clk, x, y, r, g, b);
    // KEYs are used to reset and cycle through presets
    input [3:0] KEY;
    // CLOCK_25 is used as a seed for the slower clock which controls the speed of Life generations
    input clk;
    // x and y are pixel coordinates on the 640-by-480 VGA display
    input [9:0] x, y;
    // r, g, and b represent the colour of each pixel on the VGA display
    output [3:0] r, g, b;

    /**
     * cells determines whether a square is on or off.
     * For example,
     * cells[4] == 1 means the square at the 5th column, 1st row is on.
     * cells[454] == 1 means the square at the 7th column (454 % 64 + 1 == 7), 9th row (454 / 48 == 9) is on.
     */
    wire [0:64*48-1] cells;
    // cells_reset_state and cells_preset represent the state to 
    // return all cells to when the reset KEY is pressed
    wire [0:64*48-1] cells_reset_state;
    reg [0:64*48-1] cells_preset;
    
    reg [3:0] preset_state;
    
    // This block creates presets
    initial begin
        // When the program is loaded, start with the first preset
        cells_preset[0    :64*0+63 ] <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
        cells_preset[64*1 :64*1+63 ] <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
        cells_preset[64*2 :64*2+63 ] <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
        cells_preset[64*3 :64*3+63 ] <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
        cells_preset[64*4 :64*4+63 ] <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
        cells_preset[64*5 :64*5+63 ] <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
        cells_preset[64*6 :64*6+63 ] <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
        cells_preset[64*7 :64*7+63 ] <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
        cells_preset[64*8 :64*8+63 ] <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
        cells_preset[64*9 :64*9+63 ] <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
        cells_preset[64*10:64*10+63] <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
        cells_preset[64*11:64*11+63] <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
        cells_preset[64*12:64*12+63] <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
        cells_preset[64*13:64*13+63] <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
        cells_preset[64*14:64*14+63] <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
        cells_preset[64*15:64*15+63] <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
        cells_preset[64*16:64*16+63] <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
        cells_preset[64*17:64*17+63] <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
        cells_preset[64*18:64*18+63] <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
        cells_preset[64*19:64*19+63] <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
        cells_preset[64*20:64*20+63] <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
        cells_preset[64*21:64*21+63] <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
        cells_preset[64*22:64*22+63] <= 64'b0000000000000000000000000110010000000000000000000000000000000000;
        cells_preset[64*23:64*23+63] <= 64'b0000000000000000000000000100010000000000000000000000000000000000;
        cells_preset[64*24:64*24+63] <= 64'b0000000000000000000000000100110000000000000000000000000000000000;
        cells_preset[64*25:64*25+63] <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
        cells_preset[64*26:64*26+63] <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
        cells_preset[64*27:64*27+63] <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
        cells_preset[64*28:64*28+63] <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
        cells_preset[64*29:64*29+63] <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
        cells_preset[64*30:64*30+63] <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
        cells_preset[64*31:64*31+63] <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
        cells_preset[64*32:64*32+63] <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
        cells_preset[64*33:64*33+63] <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
        cells_preset[64*34:64*34+63] <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
        cells_preset[64*35:64*35+63] <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
        cells_preset[64*36:64*36+63] <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
        cells_preset[64*37:64*37+63] <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
        cells_preset[64*38:64*38+63] <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
        cells_preset[64*39:64*39+63] <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
        cells_preset[64*40:64*40+63] <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
        cells_preset[64*41:64*41+63] <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
        cells_preset[64*42:64*42+63] <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
        cells_preset[64*43:64*43+63] <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
        cells_preset[64*44:64*44+63] <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
        cells_preset[64*45:64*45+63] <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
        cells_preset[64*46:64*46+63] <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
        cells_preset[64*47:64*47+63] <= 64'b0000000000000000000000000000000000000000000000000000000000000000;

        preset_state <= 2;
    end
    
    // When KEY[2] is pressed, cycle through presets
    /*always @(posedge KEY[2]) begin
        if (preset_state == 1) begin
            cells_preset[0    :64*0+63 ] <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
            cells_preset[64*1 :64*1+63 ] <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
            cells_preset[64*2 :64*2+63 ] <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
            cells_preset[64*3 :64*3+63 ] <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
            cells_preset[64*4 :64*4+63 ] <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
            cells_preset[64*5 :64*5+63 ] <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
            cells_preset[64*6 :64*6+63 ] <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
            cells_preset[64*7 :64*7+63 ] <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
            cells_preset[64*8 :64*8+63 ] <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
            cells_preset[64*9 :64*9+63 ] <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
            cells_preset[64*10:64*10+63] <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
            cells_preset[64*11:64*11+63] <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
            cells_preset[64*12:64*12+63] <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
            cells_preset[64*13:64*13+63] <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
            cells_preset[64*14:64*14+63] <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
            cells_preset[64*15:64*15+63] <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
            cells_preset[64*16:64*16+63] <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
            cells_preset[64*17:64*17+63] <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
            cells_preset[64*18:64*18+63] <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
            cells_preset[64*19:64*19+63] <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
            cells_preset[64*20:64*20+63] <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
            cells_preset[64*21:64*21+63] <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
            cells_preset[64*22:64*22+63] <= 64'b0000000000000000000000000110010000000000000000000000000000000000;
            cells_preset[64*23:64*23+63] <= 64'b0000000000000000000000000100010000000000000000000000000000000000;
            cells_preset[64*24:64*24+63] <= 64'b0000000000000000000000000100110000000000000000000000000000000000;
            cells_preset[64*25:64*25+63] <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
            cells_preset[64*26:64*26+63] <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
            cells_preset[64*27:64*27+63] <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
            cells_preset[64*28:64*28+63] <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
            cells_preset[64*29:64*29+63] <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
            cells_preset[64*30:64*30+63] <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
            cells_preset[64*31:64*31+63] <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
            cells_preset[64*32:64*32+63] <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
            cells_preset[64*33:64*33+63] <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
            cells_preset[64*34:64*34+63] <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
            cells_preset[64*35:64*35+63] <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
            cells_preset[64*36:64*36+63] <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
            cells_preset[64*37:64*37+63] <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
            cells_preset[64*38:64*38+63] <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
            cells_preset[64*39:64*39+63] <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
            cells_preset[64*40:64*40+63] <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
            cells_preset[64*41:64*41+63] <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
            cells_preset[64*42:64*42+63] <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
            cells_preset[64*43:64*43+63] <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
            cells_preset[64*44:64*44+63] <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
            cells_preset[64*45:64*45+63] <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
            cells_preset[64*46:64*46+63] <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
            cells_preset[64*47:64*47+63] <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
                      
            preset_state <= 2;
        end else if (preset_state == 2) begin
            cells_preset[0    :64*0+63 ] <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
            cells_preset[64*1 :64*1+63 ] <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
            cells_preset[64*2 :64*2+63 ] <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
            cells_preset[64*3 :64*3+63 ] <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
            cells_preset[64*4 :64*4+63 ] <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
            cells_preset[64*5 :64*5+63 ] <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
            cells_preset[64*6 :64*6+63 ] <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
            cells_preset[64*7 :64*7+63 ] <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
            cells_preset[64*8 :64*8+63 ] <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
            cells_preset[64*9 :64*9+63 ] <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
            cells_preset[64*10:64*10+63] <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
            cells_preset[64*11:64*11+63] <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
            cells_preset[64*12:64*12+63] <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
            cells_preset[64*13:64*13+63] <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
            cells_preset[64*14:64*14+63] <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
            cells_preset[64*15:64*15+63] <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
            cells_preset[64*16:64*16+63] <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
            cells_preset[64*17:64*17+63] <= 64'b0000000000000001100000000110000000000000000000000000000000000000;
            cells_preset[64*18:64*18+63] <= 64'b0000000000000001100000001000000000000000000000000000000000000000;
            cells_preset[64*19:64*19+63] <= 64'b0000000000000000000000000001000000000000000000000000000000000000;
            cells_preset[64*20:64*20+63] <= 64'b0000000000000000000000011010000000000000000000000000000000000000;
            cells_preset[64*21:64*21+63] <= 64'b0000000000000000000000011000000000000000000000000000000000000000;
            cells_preset[64*22:64*22+63] <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
            cells_preset[64*23:64*23+63] <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
            cells_preset[64*24:64*24+63] <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
            cells_preset[64*25:64*25+63] <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
            cells_preset[64*26:64*26+63] <= 64'b0000000000000000000000110000000000000000000000000000000000000000;
            cells_preset[64*27:64*27+63] <= 64'b0000000000000000000010110000000000000000000000000000000000000000;
            cells_preset[64*28:64*28+63] <= 64'b0000000000000000000100000000000000000000000000000000000000000000;
            cells_preset[64*29:64*29+63] <= 64'b0000000000000000000000100000001100000000000000000000000000000000;
            cells_preset[64*30:64*30+63] <= 64'b0000000000000000000011000000001100000000000000000000000000000000;
            cells_preset[64*31:64*31+63] <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
            cells_preset[64*32:64*32+63] <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
            cells_preset[64*33:64*33+63] <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
            cells_preset[64*34:64*34+63] <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
            cells_preset[64*35:64*35+63] <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
            cells_preset[64*36:64*36+63] <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
            cells_preset[64*37:64*37+63] <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
            cells_preset[64*38:64*38+63] <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
            cells_preset[64*39:64*39+63] <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
            cells_preset[64*40:64*40+63] <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
            cells_preset[64*41:64*41+63] <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
            cells_preset[64*42:64*42+63] <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
            cells_preset[64*43:64*43+63] <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
            cells_preset[64*44:64*44+63] <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
            cells_preset[64*45:64*45+63] <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
            cells_preset[64*46:64*46+63] <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
            cells_preset[64*47:64*47+63] <= 64'b0000000000000000000000000000000000000000000000000000000000000000;

            preset_state <= 3;
        end else if (preset_state == 3) begin
            cells_preset[0    :64*0+63 ] <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
            cells_preset[64*1 :64*1+63 ] <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
            cells_preset[64*2 :64*2+63 ] <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
            cells_preset[64*3 :64*3+63 ] <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
            cells_preset[64*4 :64*4+63 ] <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
            cells_preset[64*5 :64*5+63 ] <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
            cells_preset[64*6 :64*6+63 ] <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
            cells_preset[64*7 :64*7+63 ] <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
            cells_preset[64*8 :64*8+63 ] <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
            cells_preset[64*9 :64*9+63 ] <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
            cells_preset[64*10:64*10+63] <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
            cells_preset[64*11:64*11+63] <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
            cells_preset[64*12:64*12+63] <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
            cells_preset[64*13:64*13+63] <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
            cells_preset[64*14:64*14+63] <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
            cells_preset[64*15:64*15+63] <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
            cells_preset[64*16:64*16+63] <= 64'b0000000000000000000011000000110000000000000000000000000000000000;
            cells_preset[64*17:64*17+63] <= 64'b0000000000000000000100100001001000000000000000000000000000000000;
            cells_preset[64*18:64*18+63] <= 64'b0000000000000000000101000000101000000000000000000000000000000000;
            cells_preset[64*19:64*19+63] <= 64'b0000000000000000011001110011100110000000000000000000000000000000;
            cells_preset[64*20:64*20+63] <= 64'b0000000000000000100000010010000001000000000000000000000000000000;
            cells_preset[64*21:64*21+63] <= 64'b0000000000000000101100000000001101000000000000000000000000000000;
            cells_preset[64*22:64*22+63] <= 64'b0000000000000000010100000000001010000000000000000000000000000000;
            cells_preset[64*23:64*23+63] <= 64'b0000000000000000000110001100011000000000000000000000000000000000;
            cells_preset[64*24:64*24+63] <= 64'b0000000000000000000000010100000000000000000000000000000000000000;
            cells_preset[64*25:64*25+63] <= 64'b0000000000000000000000011000000000000000000000000000000000000000;
            cells_preset[64*26:64*26+63] <= 64'b0000000000000000000110000000011000000000000000000000000000000000;
            cells_preset[64*27:64*27+63] <= 64'b0000000000000000010100000000001010000000000000000000000000000000;
            cells_preset[64*28:64*28+63] <= 64'b0000000000000000101100000000001101000000000000000000000000000000;
            cells_preset[64*29:64*29+63] <= 64'b0000000000000000100000010010000001000000000000000000000000000000;
            cells_preset[64*30:64*30+63] <= 64'b0000000000000000011001110011100110000000000000000000000000000000;
            cells_preset[64*31:64*31+63] <= 64'b0000000000000000000101000000101000000000000000000000000000000000;
            cells_preset[64*32:64*32+63] <= 64'b0000000000000000000100100001001000000000000000000000000000000000;
            cells_preset[64*33:64*33+63] <= 64'b0000000000000000000011000000110000000000000000000000000000000000;
            cells_preset[64*34:64*34+63] <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
            cells_preset[64*35:64*35+63] <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
            cells_preset[64*36:64*36+63] <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
            cells_preset[64*37:64*37+63] <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
            cells_preset[64*38:64*38+63] <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
            cells_preset[64*39:64*39+63] <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
            cells_preset[64*40:64*40+63] <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
            cells_preset[64*41:64*41+63] <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
            cells_preset[64*42:64*42+63] <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
            cells_preset[64*43:64*43+63] <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
            cells_preset[64*44:64*44+63] <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
            cells_preset[64*45:64*45+63] <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
            cells_preset[64*46:64*46+63] <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
            cells_preset[64*47:64*47+63] <= 64'b0000000000000000000000000000000000000000000000000000000000000000;

            preset_state <= 4;
        end else if (preset_state == 4) begin
            cells_preset[0    :64*0+63 ] <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
            cells_preset[64*1 :64*1+63 ] <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
            cells_preset[64*2 :64*2+63 ] <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
            cells_preset[64*3 :64*3+63 ] <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
            cells_preset[64*4 :64*4+63 ] <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
            cells_preset[64*5 :64*5+63 ] <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
            cells_preset[64*6 :64*6+63 ] <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
            cells_preset[64*7 :64*7+63 ] <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
            cells_preset[64*8 :64*8+63 ] <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
            cells_preset[64*9 :64*9+63 ] <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
            cells_preset[64*10:64*10+63] <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
            cells_preset[64*11:64*11+63] <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
            cells_preset[64*12:64*12+63] <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
            cells_preset[64*13:64*13+63] <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
            cells_preset[64*14:64*14+63] <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
            cells_preset[64*15:64*15+63] <= 64'b0000000000000000000000100000000000000000000000000000000000000000;
            cells_preset[64*16:64*16+63] <= 64'b0000000000000000000001110000000000000000000000000000000000000000;
            cells_preset[64*17:64*17+63] <= 64'b0000000000000000000011010000010000000000000000000000000000000000;
            cells_preset[64*18:64*18+63] <= 64'b0000000000000000000011100000111000000000000000000000000000000000;
            cells_preset[64*19:64*19+63] <= 64'b0000000000000000000001100001001100011100000000000000000000000000;
            cells_preset[64*20:64*20+63] <= 64'b0000000000000000000000000001110000100100000000000000000000000000;
            cells_preset[64*21:64*21+63] <= 64'b0000000000000000000000000000000000000100000000000000000000000000;
            cells_preset[64*22:64*22+63] <= 64'b0000000000000000000000000000000000000100000000000000000000000000;
            cells_preset[64*23:64*23+63] <= 64'b0000000000000000000000000000000000001000000000000000000000000000;
            cells_preset[64*24:64*24+63] <= 64'b0000000000000000000001110000000000000000000000000000000000000000;
            cells_preset[64*25:64*25+63] <= 64'b0000000000000000000001001000000000000000000000000000000000000000;
            cells_preset[64*26:64*26+63] <= 64'b0000000000000000000001000000000000000000000000000000000000000000;
            cells_preset[64*27:64*27+63] <= 64'b0000000000000000000001000000000000000000000000000000000000000000;
            cells_preset[64*28:64*28+63] <= 64'b0000000000000000000000100000000000000000000000000000000000000000;
            cells_preset[64*29:64*29+63] <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
            cells_preset[64*30:64*30+63] <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
            cells_preset[64*31:64*31+63] <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
            cells_preset[64*32:64*32+63] <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
            cells_preset[64*33:64*33+63] <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
            cells_preset[64*34:64*34+63] <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
            cells_preset[64*35:64*35+63] <= 64'b0000000000000000000111000000000000000000000000000000000000000000;
            cells_preset[64*36:64*36+63] <= 64'b0000000000000000000100100000000000010000000000000000000000000000;
            cells_preset[64*37:64*37+63] <= 64'b0000000000000000000100000000000000111000000000000000000000000000;
            cells_preset[64*38:64*38+63] <= 64'b0000000000000000000100000000000001101000000000000000000000000000;
            cells_preset[64*39:64*39+63] <= 64'b0000000000000000000100000000000001110000000000000000000000000000;
            cells_preset[64*40:64*40+63] <= 64'b0000000000000000000010000000000000110000000000000000000000000000;
            cells_preset[64*41:64*41+63] <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
            cells_preset[64*42:64*42+63] <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
            cells_preset[64*43:64*43+63] <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
            cells_preset[64*44:64*44+63] <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
            cells_preset[64*45:64*45+63] <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
            cells_preset[64*46:64*46+63] <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
            cells_preset[64*47:64*47+63] <= 64'b0000000000000000000000000000000000000000000000000000000000000000;

            preset_state <= 5;
        end else if (preset_state == 5) begin
            cells_preset[0    :64*0+63 ] <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
            cells_preset[64*1 :64*1+63 ] <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
            cells_preset[64*2 :64*2+63 ] <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
            cells_preset[64*3 :64*3+63 ] <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
            cells_preset[64*4 :64*4+63 ] <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
            cells_preset[64*5 :64*5+63 ] <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
            cells_preset[64*6 :64*6+63 ] <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
            cells_preset[64*7 :64*7+63 ] <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
            cells_preset[64*8 :64*8+63 ] <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
            cells_preset[64*9 :64*9+63 ] <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
            cells_preset[64*10:64*10+63] <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
            cells_preset[64*11:64*11+63] <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
            cells_preset[64*12:64*12+63] <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
            cells_preset[64*13:64*13+63] <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
            cells_preset[64*14:64*14+63] <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
            cells_preset[64*15:64*15+63] <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
            cells_preset[64*16:64*16+63] <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
            cells_preset[64*17:64*17+63] <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
            cells_preset[64*18:64*18+63] <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
            cells_preset[64*19:64*19+63] <= 64'b0000000000110001100011000110001100011000110001100000000000000000;
            cells_preset[64*20:64*20+63] <= 64'b0000000000001100011000110001100011000110001100011000000000000000;
            cells_preset[64*21:64*21+63] <= 64'b0000000000001100011000110001100011000110001100011000000000000000;
            cells_preset[64*22:64*22+63] <= 64'b0000000000110001100011000110001100011000110001100000000000000000;
            cells_preset[64*23:64*23+63] <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
            cells_preset[64*24:64*24+63] <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
            cells_preset[64*25:64*25+63] <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
            cells_preset[64*26:64*26+63] <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
            cells_preset[64*27:64*27+63] <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
            cells_preset[64*28:64*28+63] <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
            cells_preset[64*29:64*29+63] <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
            cells_preset[64*30:64*30+63] <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
            cells_preset[64*31:64*31+63] <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
            cells_preset[64*32:64*32+63] <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
            cells_preset[64*33:64*33+63] <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
            cells_preset[64*34:64*34+63] <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
            cells_preset[64*35:64*35+63] <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
            cells_preset[64*36:64*36+63] <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
            cells_preset[64*37:64*37+63] <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
            cells_preset[64*38:64*38+63] <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
            cells_preset[64*39:64*39+63] <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
            cells_preset[64*40:64*40+63] <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
            cells_preset[64*41:64*41+63] <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
            cells_preset[64*42:64*42+63] <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
            cells_preset[64*43:64*43+63] <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
            cells_preset[64*44:64*44+63] <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
            cells_preset[64*45:64*45+63] <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
            cells_preset[64*46:64*46+63] <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
            cells_preset[64*47:64*47+63] <= 64'b0000000000000000000000000000000000000000000000000000000000000000;

            preset_state <= 1;
        end 

    end */

    // The value of cells_reset_state is the same as the current value of cells_preset
    assign cells_reset_state = cells_preset;

    // Create a clock to control the speed of generations
    //wire clk1;
    //clk_div(.clk(clk), .q(clk1));
    //wire enable;
    wire use_enable;
    
    clk_div div(.clk(clk), .en(use_enable));
    //dff_en dff_en(.DFF_CLK(clk), .clock_en(enable), .Q(use_enable));
    
    /**
     * Assign neighbours for each cell depending on the cell's location.
     * Cells on the edges and corners of the grid must be dealt with separately since
     * their neighbours are not directly adjacent.
     */
    genvar i;
    generate
        for (i = 0; i < 64 * 48; i = i + 1) begin : CELLS
            wire [7:0] neighbours;
            if (i == 0) begin
                // Top-left square
                assign neighbours[0] = cells[64*48 - 1];
                assign neighbours[1] = cells[64*48 - 64];
                assign neighbours[2] = cells[64*48 - 64 + 1];
                assign neighbours[3] = cells[i     + 64 - 1];
                assign neighbours[4] = cells[i     + 1];
                assign neighbours[5] = cells[64    + 64 - 1];
                assign neighbours[6] = cells[64];
                assign neighbours[7] = cells[64    + 1];
            end else if (i == 63) begin
                // Top-right square
                assign neighbours[0] = cells[64*48 - 1 - 1];
                assign neighbours[1] = cells[64*48 - 1];
                assign neighbours[2] = cells[64*48 - 64];
                assign neighbours[3] = cells[i     - 1];
                assign neighbours[4] = cells[0];
                assign neighbours[5] = cells[i     + 64 - 1];
                assign neighbours[6] = cells[i     + 64];
                assign neighbours[7] = cells[i     + 1];
            end else if (i == 64*48 - 64) begin
                // Bottom-left square
                assign neighbours[0] = cells[i - 1];
                assign neighbours[1] = cells[i - 64];
                assign neighbours[2] = cells[i - 64 + 1];
                assign neighbours[3] = cells[i + 64 - 1];
                assign neighbours[4] = cells[i + 1];
                assign neighbours[5] = cells[0 + 64 - 1];
                assign neighbours[6] = cells[0];
                assign neighbours[7] = cells[0 + 1];
            end else if (i == 64*48 - 1) begin
                // Bottom-right square
                assign neighbours[0] = cells[i - 64 - 1];
                assign neighbours[1] = cells[i - 64];
                assign neighbours[2] = cells[i - 64 - 64 + 1];
                assign neighbours[3] = cells[i - 1];
                assign neighbours[4] = cells[i - 64 + 1];
                assign neighbours[5] = cells[0 + 64 - 1 - 1];
                assign neighbours[6] = cells[0 + 64 - 1];
                assign neighbours[7] = cells[0];
            end else if (i < 63) begin
                // Top row
                assign neighbours[0] = cells[64*48 - 64 + i - 1];
                assign neighbours[1] = cells[64*48 - 64 + i];
                assign neighbours[2] = cells[64*48 - 64 + i + 1];
                assign neighbours[3] = cells[i - 1];
                assign neighbours[4] = cells[i + 1];
                assign neighbours[5] = cells[i + 64 - 1];
                assign neighbours[6] = cells[i + 64];
                assign neighbours[7] = cells[i + 64 + 1];
            end else if (i > 64*48 - 64) begin
                // Bottom row
                assign neighbours[0] = cells[i - 64 - 1];
                assign neighbours[1] = cells[i - 64];
                assign neighbours[2] = cells[i - 64 + 1];
                assign neighbours[3] = cells[i - 1];
                assign neighbours[4] = cells[i + 1];
                assign neighbours[5] = cells[0 + i - 1];
                assign neighbours[6] = cells[0 + i];
                assign neighbours[7] = cells[0 + i + 1];
            end else if (i % 64 == 0) begin
                // Leftmost column
                assign neighbours[0] = cells[i - 1];
                assign neighbours[1] = cells[i - 64];
                assign neighbours[2] = cells[i - 64 + 1];
                assign neighbours[3] = cells[i + 64 - 1];
                assign neighbours[4] = cells[i + 1];
                assign neighbours[5] = cells[i + 64 + 64 - 1];
                assign neighbours[6] = cells[i + 64];
                assign neighbours[7] = cells[i + 64 + 1];
            end else if ((i + 1) % 64 == 0) begin
                // Rightmost column
                assign neighbours[0] = cells[i - 64 - 1];
                assign neighbours[1] = cells[i - 64];
                assign neighbours[2] = cells[i - 64 - 64 + 1];
                assign neighbours[3] = cells[i - 1];
                assign neighbours[4] = cells[i - 64 + 1];
                assign neighbours[5] = cells[i + 64 - 1];
                assign neighbours[6] = cells[i + 64];
                assign neighbours[7] = cells[i + 1];
            end else begin
                // Middle squares
                assign neighbours[0] = cells[i - 64 - 1];
                assign neighbours[1] = cells[i - 64];
                assign neighbours[2] = cells[i - 64 + 1];
                assign neighbours[3] = cells[i - 1];
                assign neighbours[4] = cells[i + 1];
                assign neighbours[5] = cells[i + 64 - 1];
                assign neighbours[6] = cells[i + 64];
                assign neighbours[7] = cells[i + 64 + 1];
            end
            // Create the module for the cell
            live_cell(.neighbours(neighbours), .clk(clk), .use_enable(use_enable), .Rst(KEY[2]), .initial_state(cells_reset_state[i]), .state(cells[i]));
        end
    endgenerate
        
    // Show the cells on the VGA display
    display_grid(.cells(cells), .x(x), .y(y), .r(r), .g(g), .b(b));

endmodule